(** * Natural Transformations *)
(** Since there are only notations in [NaturalTransformation.Notations], we can just export those. *)
Require Export NaturalTransformation.Notations.

(** ** Definition of natural transformation *)
Require NaturalTransformation.Core.
(** ** Composition of natural transformations *)
Require NaturalTransformation.Composition.Core.
(** ** Dual natural transformations *)
Require NaturalTransformation.Dual.
(** ** Identity natural transformation *)
Require NaturalTransformation.Identity.
(** ** Natural isomorphisms *)
Require NaturalTransformation.Isomorphisms.
(** ** Path space of natural transformation type *)
Require NaturalTransformation.Paths.
(** ** Pointwise natural transformations *)
Require NaturalTransformation.Pointwise.
(** ** Sums of natural transformations *)
Require NaturalTransformation.Sum.
(** ** Products of natural transformations *)
Require NaturalTransformation.Prod.

Include NaturalTransformation.Core.
Include NaturalTransformation.Composition.Core.
Include NaturalTransformation.Dual.
Include NaturalTransformation.Identity.
Include NaturalTransformation.Isomorphisms.
Include NaturalTransformation.Paths.
Include NaturalTransformation.Pointwise.
Include NaturalTransformation.Sum.
Include NaturalTransformation.Prod.
(** We don't want to make utf-8 notations the default, so we don't export them. *)

(** Since [Composition] is a separate sub-directory, we need to re-create the module structure *)
Module Composition.
  Require NaturalTransformation.Composition.Composition.
  Include NaturalTransformation.Composition.Composition.
End Composition.
